// LUT for the big boi
module loot
(
  output cs,
  output modes,

  input clk
);
endmodule

// LUT for the smoller baby
module lute
(
  input cs,
  input clk
);
endmodule
