`include "datamemory.v"
`include "dflipflop.v"
`include "inputconditioner.v"
`include "LUT.v"

module baby(
  input miso,
  input address,
  output mosi,
  output sclk,
  output cs
);
 wire 



shiftregister8 schwifty ();
