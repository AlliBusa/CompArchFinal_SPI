// LUT for
module loot
(
  output cs,
  output modes,

  input clk
);
endmodule

module lute
(
  input cs,
  input clk
);
endmodule
